module animals

import core

pub struct Funny {
	id             int
	genes          core.GeneSequence
	generation_nbr int
}
