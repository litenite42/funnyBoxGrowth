module interfaces

pub interface IEntity {
	id int
}
